-------------------------------------------------------------------------------
-- MEL Counter Project - Top Level Testbench Entity                         --
--                                                                           --
-- Description: Testbench entity for the complete counter system            --
--              verification. Tests integration of IO control and           --
--              counter units with realistic switch scenarios.              --
--                                                                           --
-- Author : Summer Paulus, Matthias Brinskelle                              --
-- Date : 18.06.2025                                                        --
-- File : tb_cntr_top_.vhd                                                  --
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_cntr_top is
  -- Testbench has no ports
end tb_cntr_top;
