-------------------------------------------------------------------------------
-- MEL Counter Project - Counter Unit Testbench Entity                      --
--                                                                           --
-- Description: Testbench entity for the counter unit verification.         --
--              Tests counting functionality, priority control, and          --
--              wraparound behavior for octal counter.                      --
--                                                                           --
-- Author : Summer Paulus, Matthias Brinskelle                              --
-- Date : 18.06.2025                                                        --
-- File : tb_cntr_.vhd                                                      --
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_cntr is
  -- Testbench has no ports
end tb_cntr;
