-------------------------------------------------------------------------------
-- MEL Counter Project - Counter Unit Configuration                         --
--                                                                           --
-- Description: Configuration file binding the cntr entity to its           --
--              RTL architecture implementation.                            --
--                                                                           --
-- Author : Summer Paulus, Matthias Brinskelle                              --
-- Date : 18.06.2025                                                        --
-- File : cntr_rtl_cfg.vhd                                                 --
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

configuration cntr_rtl_cfg of cntr is
  for rtl
  end for;
end cntr_rtl_cfg;
