-------------------------------------------------------------------------------
-- MEL Counter Project - IO Control Unit Testbench Entity                   --
--                                                                           --
-- Description: Testbench entity for the IO control unit verification.      --
--              Tests debouncing, 7-segment display, and LED functionality.  --
--                                                                           --
-- Author : Summer Paulus, Matthias Brinskelle                              --
-- Date : 18.06.2025                                                        --
-- File : tb_io_ctrl_.vhd                                                   --
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity tb_io_ctrl is
  -- Testbench has no ports
end tb_io_ctrl;
