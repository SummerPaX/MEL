-------------------------------------------------------------------------------
-- VHDL Class Example Fulladder, Design                                      --
--                                                                           --
-- Description: This is the configuration for the entity orgate and the      --
--              architecture rtl.                                            --
--                                                                           --
-- Author : Paulus Summer, Matthias Brinskelle                               --
-- Date : 18.06.2025                                                         --
-- File : orgate_rtl_cfg.vhd                                                 --
-------------------------------------------------------------------------------

configuration orgate_rtl_cfg of orgate is
  for rtl  -- architecture rtl is used for entity orgate
  end for;
end orgate_rtl_cfg;
