-------------------------------------------------------------------------------
-- MEL Counter Project - IO Control Unit Testbench Entity                    --
--                                                                           --
-- Description: Testbench entity for the IO control unit verification.       --
--              Tests debouncing, 7-segment display, and LED functionality.  --
--                                                                           --
-- Author : Summer Paulus, Matthias Brinskelle                               --
-- Date : 19.06.2025                                                         --
-- File : tb_io_ctrl_.vhd                                                    --
-------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY tb_io_ctrl IS
END tb_io_ctrl;