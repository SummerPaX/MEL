-------------------------------------------------------------------------------
-- MEL Counter Project - Top Level Testbench Entity                          --
--                                                                           --
-- Description: Testbench entity for the complete counter system             --
--              verification. Tests integration of IO control and            --
--              counter units with realistic switch scenarios.               --
--                                                                           --
-- Author : Summer Paulus, Matthias Brinskelle                               --
-- Date : 19.06.2025                                                         --
-- File : tb_cntr_top_.vhd                                                   --
-------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY tb_cntr_top IS
END tb_cntr_top;