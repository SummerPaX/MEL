-------------------------------------------------------------------------------
-- VHDL Class Example Fulladder, Design                                      --
--                                                                           --
-- Description: This is the configuration for the entity halfadder and the   --
--              architecture rtl.                                            --
--                                                                           --
-- Author : Paulus Summer, Matthias Brinskelle                               --
-- Date : 18.06.2025                                                         --
-- File : halfadder_rtl_cfg.vhd                                              --
-------------------------------------------------------------------------------

configuration halfadder_rtl_cfg of halfadder is
  for rtl  -- architecture rtl is used for entity halfadder
  end for;
end halfadder_rtl_cfg;
