-------------------------------------------------------------------------------
-- VHDL Class Example Fulladder, Design                                      --
--                                                                           --
-- Description: This is the configuration for the entity fulladder and the   --
--              architecture struc.                                          --
--                                                                           --
-- Author : Paulus Summer, Matthias Brinskelle                               --
-- Date : 18.06.2025                                                         --
-- File : fulladder_struc_cfg.vhd                                            --
-------------------------------------------------------------------------------

configuration fulladder_struc_cfg of fulladder is
  for struc -- architecture struc is used for entity fulladder
  end for;
end fulladder_struc_cfg;
