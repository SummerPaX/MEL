-------------------------------------------------------------------------------
-- MEL Counter Project - Counter Unit Testbench Entity                       --
--                                                                           --
-- Description: Testbench entity declaration for the counter unit.           --
--              Tests all counter functionality including up/down counting,  --
--              clear, hold, and wraparound behavior.                        --
--                                                                           --
-- Author : Summer Paulus, Matthias Brinskelle                               --
-- Date : 19.06.2025                                                         --
-- File : tb_cntr_.vhd                                                       --
-------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY tb_cntr IS
  -- Testbench has no ports
END tb_cntr;